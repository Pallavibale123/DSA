module testbench;
  //automatic makes Each call gets its own copy of local variables. Local variables are stack-allocated and disappear when the function call ends
  function automatic int count_setbits(input int unsigned n);

    int count = 0;
    while (n != 0)begin
      n = n & (n-1);
      count = count + 1;
    end
    return count;
    
  endfunction
  
  initial begin
    int unsigned num;
    int result;
	int unsigned testing[7:0] = '{32'd0, 32'd1, 32'd2, 32'hFFFFFFFF, 32'd7, 32'd64, 32'd16, 32'd15};
    
    foreach (testing[i])begin
      num = testing[i];
      result = count_setbits(num);
      $display("The total number of 1's is = %0d for number = %0d", result, num);
    end
    $finish;
  end
  
endmodule

/*
The total number of 1's is = 0 for number = 0
The total number of 1's is = 1 for number = 1
The total number of 1's is = 1 for number = 2
The total number of 1's is = 32 for number = 4294967295
The total number of 1's is = 3 for number = 7
The total number of 1's is = 1 for number = 64
The total number of 1's is = 1 for number = 16
The total number of 1's is = 4 for number = 15
*/
